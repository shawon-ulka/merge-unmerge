Hello
this is an spice file

.start


.end